magic
tech sky130A
magscale 1 2
timestamp 1756664610
<< isosubstrate >>
rect 2174 -8984 2178 -7880
rect 2174 -8992 3156 -8984
<< nwell >>
rect 3680 -7910 3708 -7900
rect 3578 -7976 3708 -7910
rect 3794 -7970 3860 -7824
rect 3418 -8206 3504 -8000
rect 3638 -8244 3708 -7976
rect 2854 -8258 2864 -8246
rect 3578 -8302 3708 -8244
rect 3578 -8308 3680 -8302
rect 3576 -8328 4108 -8308
rect 3576 -8376 3894 -8328
<< pwell >>
rect 3294 -8462 3310 -8458
rect 2422 -8540 2430 -8482
rect 2440 -8664 2468 -8516
rect 2472 -8634 2538 -8580
rect 2580 -8634 2646 -8580
rect 2440 -8682 2474 -8664
rect 2854 -8670 2902 -8494
rect 3002 -8634 3146 -8568
rect 3294 -8592 3312 -8462
rect 3292 -8644 3312 -8592
rect 3470 -8620 3536 -8562
rect 3920 -8628 3940 -8470
rect 3292 -8650 3376 -8644
rect 3624 -8650 3706 -8634
rect 3064 -8754 3134 -8678
rect 3292 -8740 3482 -8650
rect 3624 -8662 3796 -8650
rect 2580 -8854 2646 -8788
rect 3312 -8838 3476 -8740
rect 3312 -8866 3376 -8838
rect 3530 -8842 3796 -8662
rect 3624 -8844 3796 -8842
rect 3624 -8860 3746 -8844
rect 3920 -8846 3934 -8628
rect 3952 -8662 4006 -8646
rect 3952 -8844 4108 -8662
rect 3952 -8856 4008 -8844
rect 4162 -8850 4328 -8654
rect 4958 -8862 5106 -8660
rect 3468 -8940 4168 -8878
rect 3404 -8982 3596 -8968
rect 3288 -9038 4322 -8982
rect 4696 -9038 4706 -8994
rect 4846 -9002 4872 -8986
rect 5072 -9002 5142 -8970
rect 4846 -9008 5010 -9002
rect 4846 -9038 4872 -9008
rect 3288 -9108 5046 -9038
rect 3288 -9174 4322 -9108
<< psubdiff >>
rect 4852 -9008 5010 -9002
<< poly >>
rect 2376 -8312 2520 -8240
rect 2910 -8246 2940 -8208
rect 2794 -8302 2940 -8246
rect 2472 -8634 2538 -8580
rect 2440 -8856 2520 -8790
rect 2796 -8858 2940 -8792
<< locali >>
rect 4436 -8072 4472 -7918
rect 3070 -8642 3104 -8590
rect 3070 -8846 3104 -8748
rect 3328 -8838 3362 -8660
rect 3642 -8662 3680 -8648
rect 3960 -8838 3994 -8662
rect 4442 -8672 4474 -8584
rect 4442 -8940 4474 -8858
rect 3422 -9000 3424 -8990
rect 3898 -9000 3900 -8990
rect 4054 -9000 4056 -8992
rect 5072 -9000 5106 -8970
<< viali >>
rect 3532 -7858 3690 -7824
rect 3848 -7858 4006 -7824
rect 4534 -7856 4692 -7822
rect 4848 -7856 5008 -7820
rect 2432 -7966 2484 -7932
rect 2848 -7966 2908 -7932
rect 3436 -8196 3472 -8018
rect 3752 -8196 3786 -8018
rect 4436 -8290 4472 -8072
rect 4754 -8186 4788 -8028
rect 2430 -8528 2482 -8494
rect 2852 -8528 2904 -8494
rect 3070 -8742 3104 -8658
rect 3642 -8824 3680 -8662
rect 4276 -8838 4310 -8662
rect 4442 -8858 4476 -8672
rect 4758 -8850 4792 -8684
rect 3424 -9024 3582 -8990
rect 3740 -9024 3898 -8990
rect 4056 -9024 4214 -8990
rect 4536 -9036 4694 -9002
rect 4852 -9036 5010 -9002
rect 5228 -9154 5398 -8988
<< metal1 >>
rect 3118 -7720 3318 -7636
rect 2930 -7722 3318 -7720
rect 3926 -7722 4074 -7718
rect 4518 -7722 5018 -7720
rect 2930 -7780 5018 -7722
rect 2930 -7892 3020 -7780
rect 3118 -7836 3318 -7780
rect 3518 -7824 3702 -7780
rect 3770 -7782 5018 -7780
rect 3518 -7858 3532 -7824
rect 3690 -7858 3702 -7824
rect 3518 -7874 3702 -7858
rect 3820 -7824 4074 -7782
rect 4140 -7784 5018 -7782
rect 4140 -7788 4704 -7784
rect 3820 -7858 3848 -7824
rect 4006 -7858 4074 -7824
rect 3820 -7874 4074 -7858
rect 4518 -7822 4704 -7788
rect 4518 -7856 4534 -7822
rect 4692 -7856 4704 -7822
rect 4518 -7872 4704 -7856
rect 4840 -7820 5018 -7784
rect 4840 -7856 4848 -7820
rect 5008 -7856 5018 -7820
rect 5154 -7770 5354 -7652
rect 5154 -7830 5174 -7770
rect 5236 -7772 5354 -7770
rect 5236 -7830 5276 -7772
rect 5154 -7832 5276 -7830
rect 5338 -7832 5354 -7772
rect 5154 -7852 5354 -7832
rect 4840 -7872 5018 -7856
rect 2424 -7922 2494 -7920
rect 2424 -7974 2430 -7922
rect 2486 -7974 2494 -7922
rect 2424 -7978 2494 -7974
rect 2836 -7924 3020 -7892
rect 4352 -7910 4646 -7908
rect 2836 -7976 2848 -7924
rect 2908 -7976 3020 -7924
rect 3578 -7976 3684 -7910
rect 3882 -7970 3970 -7910
rect 3894 -7976 3960 -7970
rect 4190 -7974 4646 -7910
rect 4896 -7974 4960 -7908
rect 4190 -7976 4238 -7974
rect 4426 -7976 4488 -7974
rect 2836 -7978 3020 -7976
rect 3418 -8018 3592 -8004
rect 2472 -8026 2538 -8018
rect 2472 -8074 2958 -8026
rect 2424 -8120 2490 -8112
rect 2294 -8256 2344 -8128
rect 2424 -8208 2432 -8120
rect 2484 -8208 2490 -8120
rect 2752 -8126 2798 -8116
rect 2424 -8218 2490 -8208
rect 2534 -8218 2570 -8126
rect 2720 -8216 2798 -8126
rect 2844 -8122 2910 -8114
rect 2844 -8210 2850 -8122
rect 2902 -8210 2910 -8122
rect 2844 -8216 2910 -8210
rect 2954 -8126 2990 -8114
rect 2954 -8216 3040 -8126
rect 3418 -8196 3436 -8018
rect 3472 -8196 3592 -8018
rect 3418 -8206 3592 -8196
rect 2294 -8302 2520 -8256
rect 2294 -8422 2344 -8302
rect 2720 -8420 2764 -8216
rect 2794 -8302 2864 -8246
rect 2990 -8382 3040 -8216
rect 3638 -8208 3684 -7976
rect 3732 -8018 3902 -8008
rect 3732 -8196 3752 -8018
rect 3786 -8196 3902 -8018
rect 4190 -8020 4236 -7976
rect 3638 -8238 3680 -8208
rect 3732 -8210 3902 -8196
rect 3952 -8200 4236 -8020
rect 3578 -8250 3680 -8238
rect 3894 -8246 3960 -8238
rect 3568 -8314 3578 -8250
rect 3662 -8254 3680 -8250
rect 3662 -8304 3678 -8254
rect 3710 -8304 3960 -8246
rect 3662 -8314 3672 -8304
rect 3710 -8378 3756 -8304
rect 3430 -8380 3756 -8378
rect 3142 -8382 3756 -8380
rect 2990 -8392 3756 -8382
rect 4190 -8342 4236 -8200
rect 4426 -8070 4492 -8060
rect 4534 -8070 4592 -8006
rect 4426 -8072 4592 -8070
rect 4426 -8290 4436 -8072
rect 4472 -8208 4592 -8072
rect 4640 -8206 4720 -8002
rect 4750 -8020 4908 -8010
rect 4748 -8028 4908 -8020
rect 4748 -8186 4754 -8028
rect 4788 -8186 4908 -8028
rect 4748 -8192 4908 -8186
rect 4944 -8192 4954 -8016
rect 5008 -8192 5018 -8016
rect 4750 -8202 4908 -8192
rect 4472 -8290 4484 -8208
rect 4686 -8236 4720 -8206
rect 4686 -8240 4962 -8236
rect 4426 -8306 4484 -8290
rect 4582 -8342 4646 -8246
rect 2990 -8420 3758 -8392
rect 2294 -8454 2602 -8422
rect 2720 -8432 3758 -8420
rect 4190 -8400 4646 -8342
rect 4686 -8302 4964 -8240
rect 4686 -8346 4766 -8302
rect 4190 -8432 4236 -8400
rect 2720 -8434 3286 -8432
rect 2720 -8448 3028 -8434
rect 2294 -8680 2344 -8454
rect 2420 -8484 2490 -8482
rect 2420 -8536 2428 -8484
rect 2484 -8536 2490 -8484
rect 2420 -8540 2490 -8536
rect 2472 -8634 2538 -8580
rect 2424 -8674 2490 -8668
rect 2294 -8756 2378 -8680
rect 2424 -8762 2430 -8674
rect 2482 -8762 2490 -8674
rect 2570 -8680 2602 -8454
rect 2536 -8756 2602 -8680
rect 2730 -8454 3028 -8448
rect 2730 -8680 2762 -8454
rect 2842 -8484 2914 -8482
rect 2842 -8536 2850 -8484
rect 2906 -8536 2914 -8484
rect 2842 -8540 2914 -8536
rect 2892 -8640 2954 -8584
rect 2990 -8664 3028 -8454
rect 3884 -8464 4236 -8432
rect 3470 -8620 3536 -8562
rect 3786 -8620 3852 -8562
rect 2844 -8674 2910 -8668
rect 2730 -8756 2798 -8680
rect 2424 -8768 2490 -8762
rect 2844 -8762 2850 -8674
rect 2902 -8762 2910 -8674
rect 2980 -8680 3028 -8664
rect 2956 -8694 2986 -8680
rect 2990 -8758 3028 -8680
rect 3064 -8652 3110 -8646
rect 3884 -8650 3940 -8464
rect 4102 -8620 4168 -8562
rect 4582 -8576 4646 -8400
rect 4724 -8544 4766 -8346
rect 4688 -8574 4766 -8544
rect 4582 -8632 4650 -8576
rect 4688 -8632 4964 -8574
rect 4688 -8634 4924 -8632
rect 4688 -8636 4766 -8634
rect 3258 -8652 3482 -8650
rect 3064 -8658 3482 -8652
rect 3064 -8742 3070 -8658
rect 3104 -8740 3482 -8658
rect 3626 -8662 3796 -8650
rect 3874 -8652 3940 -8650
rect 3104 -8742 3110 -8740
rect 3064 -8754 3110 -8742
rect 2844 -8768 2910 -8762
rect 2376 -8976 2442 -8800
rect 2796 -8892 2862 -8802
rect 3430 -8838 3476 -8740
rect 3530 -8824 3642 -8662
rect 3680 -8824 3796 -8662
rect 3530 -8842 3796 -8824
rect 3746 -8844 3796 -8842
rect 3844 -8846 3940 -8652
rect 3876 -8848 3940 -8846
rect 3980 -8662 4086 -8648
rect 4162 -8662 4328 -8654
rect 3980 -8680 4108 -8662
rect 3980 -8820 4052 -8680
rect 4108 -8820 4118 -8680
rect 3980 -8844 4108 -8820
rect 4162 -8838 4276 -8662
rect 4310 -8838 4328 -8662
rect 3980 -8850 4096 -8844
rect 4162 -8850 4328 -8838
rect 4432 -8672 4488 -8656
rect 4688 -8662 4722 -8636
rect 3980 -8878 4050 -8850
rect 4432 -8858 4442 -8672
rect 4476 -8674 4488 -8672
rect 4676 -8674 4720 -8662
rect 4476 -8856 4590 -8674
rect 4642 -8850 4720 -8674
rect 4750 -8684 4910 -8670
rect 4750 -8850 4758 -8684
rect 4792 -8850 4910 -8684
rect 4948 -8850 4958 -8674
rect 5012 -8850 5022 -8674
rect 4476 -8858 4488 -8856
rect 2794 -8976 2864 -8892
rect 3468 -8940 4168 -8878
rect 4432 -8882 4488 -8858
rect 4750 -8862 4910 -8850
rect 4582 -8946 4650 -8890
rect 4896 -8948 4964 -8892
rect 2312 -9176 2512 -8976
rect 2730 -9176 2930 -8976
rect 5212 -8982 5600 -8970
rect 3288 -8990 4322 -8982
rect 3288 -9024 3424 -8990
rect 3582 -9024 3740 -8990
rect 3898 -9024 4056 -8990
rect 4214 -9000 4322 -8990
rect 5212 -8988 5474 -8982
rect 4530 -9000 4700 -8996
rect 4844 -9000 5018 -8996
rect 5212 -9000 5228 -8988
rect 4214 -9002 5228 -9000
rect 4214 -9024 4536 -9002
rect 3288 -9036 4536 -9024
rect 4694 -9036 4852 -9002
rect 5010 -9036 5228 -9002
rect 3288 -9154 5228 -9036
rect 5398 -9052 5474 -8988
rect 5566 -9052 5600 -8982
rect 5398 -9090 5600 -9052
rect 5398 -9154 5474 -9090
rect 3288 -9164 5474 -9154
rect 5566 -9164 5600 -9090
rect 3288 -9170 5600 -9164
rect 3288 -9174 4322 -9170
<< via1 >>
rect 5174 -7830 5236 -7770
rect 5276 -7832 5338 -7772
rect 2430 -7932 2486 -7922
rect 2430 -7966 2432 -7932
rect 2432 -7966 2484 -7932
rect 2484 -7966 2486 -7932
rect 2430 -7974 2486 -7966
rect 2848 -7932 2908 -7924
rect 2848 -7966 2908 -7932
rect 2848 -7976 2908 -7966
rect 2432 -8208 2484 -8120
rect 2850 -8210 2902 -8122
rect 3578 -8314 3662 -8250
rect 4954 -8192 5008 -8016
rect 2428 -8494 2484 -8484
rect 2428 -8528 2430 -8494
rect 2430 -8528 2482 -8494
rect 2482 -8528 2484 -8494
rect 2428 -8536 2484 -8528
rect 2430 -8762 2482 -8674
rect 2850 -8494 2906 -8484
rect 2850 -8528 2852 -8494
rect 2852 -8528 2904 -8494
rect 2904 -8528 2906 -8494
rect 2850 -8536 2906 -8528
rect 2850 -8762 2902 -8674
rect 4052 -8820 4108 -8680
rect 4958 -8850 5012 -8674
rect 5474 -9052 5566 -8982
rect 5474 -9164 5566 -9090
<< metal2 >>
rect 5156 -7770 5356 -7746
rect 5156 -7830 5174 -7770
rect 5236 -7830 5274 -7770
rect 5336 -7772 5356 -7770
rect 5156 -7832 5276 -7830
rect 5338 -7832 5356 -7772
rect 5156 -7850 5356 -7832
rect 2424 -7922 2494 -7920
rect 2424 -7974 2430 -7922
rect 2486 -7974 2494 -7922
rect 2424 -7978 2494 -7974
rect 2836 -7924 2920 -7914
rect 2836 -7976 2848 -7924
rect 2908 -7976 2920 -7924
rect 2440 -8112 2476 -7978
rect 2836 -7986 2920 -7976
rect 2424 -8120 2490 -8112
rect 2860 -8114 2894 -7986
rect 4950 -8004 5006 -7996
rect 4950 -8006 5008 -8004
rect 5006 -8016 5018 -8006
rect 2424 -8208 2432 -8120
rect 2484 -8208 2490 -8120
rect 2424 -8218 2490 -8208
rect 2844 -8122 2910 -8114
rect 2844 -8210 2850 -8122
rect 2902 -8210 2910 -8122
rect 2844 -8216 2910 -8210
rect 5008 -8192 5018 -8016
rect 5006 -8206 5018 -8192
rect 4950 -8216 5006 -8206
rect 3578 -8250 3662 -8240
rect 3576 -8314 3578 -8308
rect 3662 -8314 3680 -8250
rect 3576 -8338 3680 -8314
rect 3576 -8374 4108 -8338
rect 3576 -8376 3894 -8374
rect 2422 -8484 2490 -8482
rect 2422 -8536 2428 -8484
rect 2484 -8536 2490 -8484
rect 2422 -8540 2490 -8536
rect 2842 -8484 2914 -8482
rect 2842 -8536 2850 -8484
rect 2906 -8536 2914 -8484
rect 2842 -8540 2914 -8536
rect 2430 -8668 2482 -8540
rect 2854 -8668 2902 -8540
rect 2426 -8674 2488 -8668
rect 2426 -8762 2430 -8674
rect 2482 -8762 2488 -8674
rect 2426 -8768 2488 -8762
rect 2844 -8674 2910 -8668
rect 2844 -8762 2850 -8674
rect 2902 -8762 2910 -8674
rect 4050 -8680 4108 -8374
rect 4958 -8660 5014 -8650
rect 4050 -8752 4052 -8680
rect 2844 -8768 2910 -8762
rect 4052 -8830 4108 -8820
rect 4956 -8850 4958 -8674
rect 5014 -8850 5020 -8674
rect 4958 -8870 5014 -8860
rect 5450 -8982 5586 -8970
rect 5450 -9052 5474 -8982
rect 5566 -9052 5586 -8982
rect 5450 -9090 5586 -9052
rect 5450 -9164 5474 -9090
rect 5566 -9164 5586 -9090
rect 5450 -9170 5586 -9164
<< via2 >>
rect 5174 -7830 5236 -7770
rect 5274 -7772 5336 -7770
rect 5274 -7830 5276 -7772
rect 5276 -7830 5336 -7772
rect 4950 -8016 5006 -8006
rect 4950 -8192 4954 -8016
rect 4954 -8192 5006 -8016
rect 4950 -8206 5006 -8192
rect 4958 -8674 5014 -8660
rect 4958 -8850 5012 -8674
rect 5012 -8850 5014 -8674
rect 4958 -8860 5014 -8850
rect 5474 -9052 5566 -8982
rect 5474 -9164 5566 -9090
<< metal3 >>
rect 5156 -7766 5356 -7746
rect 5156 -7836 5168 -7766
rect 5238 -7836 5272 -7766
rect 5342 -7836 5356 -7766
rect 5156 -7852 5356 -7836
rect 4940 -8006 5016 -8001
rect 4940 -8206 4950 -8006
rect 5006 -8010 5016 -8006
rect 5016 -8198 5026 -8010
rect 5006 -8206 5016 -8198
rect 4940 -8211 5016 -8206
rect 4946 -8864 4956 -8652
rect 5022 -8864 5032 -8652
rect 4948 -8865 5024 -8864
rect 5450 -8982 5586 -8970
rect 5450 -9052 5474 -8982
rect 5566 -9052 5586 -8982
rect 5450 -9090 5586 -9052
rect 5450 -9164 5474 -9090
rect 5566 -9164 5586 -9090
rect 5450 -9172 5586 -9164
<< via3 >>
rect 5168 -7770 5238 -7766
rect 5168 -7830 5174 -7770
rect 5174 -7830 5236 -7770
rect 5236 -7830 5238 -7770
rect 5168 -7836 5238 -7830
rect 5272 -7770 5342 -7766
rect 5272 -7830 5274 -7770
rect 5274 -7830 5336 -7770
rect 5336 -7830 5342 -7770
rect 5272 -7836 5342 -7830
rect 4950 -8198 5006 -8010
rect 5006 -8198 5016 -8010
rect 4956 -8660 5022 -8652
rect 4956 -8860 4958 -8660
rect 4958 -8860 5014 -8660
rect 5014 -8860 5022 -8660
rect 4956 -8864 5022 -8860
rect 5474 -9052 5566 -8982
rect 5474 -9164 5566 -9090
<< metal4 >>
rect 5154 -7766 5356 -7746
rect 5154 -7836 5168 -7766
rect 5238 -7836 5272 -7766
rect 5342 -7836 5356 -7766
rect 5154 -7968 5356 -7836
rect 4948 -8008 5010 -7994
rect 5154 -8008 5354 -7968
rect 4948 -8010 5310 -8008
rect 4948 -8198 4950 -8010
rect 5016 -8196 5310 -8010
rect 5016 -8198 5017 -8196
rect 4948 -8199 5017 -8198
rect 4948 -8210 5010 -8199
rect 5132 -8202 5310 -8196
rect 5160 -8208 5310 -8202
rect 5246 -8240 5310 -8208
rect 4955 -8652 5023 -8651
rect 5220 -8652 5320 -8452
rect 4955 -8864 4956 -8652
rect 5022 -8864 5320 -8652
rect 4955 -8865 5023 -8864
rect 5228 -8866 5320 -8864
rect 5592 -8970 5792 -8472
rect 5450 -8982 5792 -8970
rect 5450 -9052 5474 -8982
rect 5566 -9052 5792 -8982
rect 5450 -9090 5792 -9052
rect 5450 -9164 5474 -9090
rect 5566 -9164 5792 -9090
rect 5450 -9170 5792 -9164
rect 5592 -9172 5792 -9170
use sky130_fd_pr__cap_mim_m3_1_9482M8  XC8
timestamp 1755446217
transform -1 0 5906 0 -1 -8334
box -686 -240 686 240
use sky130_fd_pr__nfet_01v8_TGNW9T  XM1
timestamp 1755446217
transform 1 0 4135 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_3SNH8H  XM2
timestamp 1755446217
transform 1 0 2877 0 1 -8718
box -263 -260 263 260
use sky130_fd_pr__pfet_01v8_J8PPQP  XM3
timestamp 1755446217
transform 1 0 3611 0 1 -8107
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_J8PPQP  XM4
timestamp 1755446217
transform 1 0 4613 0 1 -8105
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_TGNW9T  XM5
timestamp 1755446217
transform 1 0 3503 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_X8MKUN  XM6
timestamp 1755446217
transform 1 0 2877 0 1 -8165
box -263 -269 263 269
use sky130_fd_pr__nfet_01v8_TGNW9T  XM7
timestamp 1755446217
transform 1 0 3819 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_3SNH8H  XM8
timestamp 1755446217
transform 1 0 2457 0 1 -8718
box -263 -260 263 260
use sky130_fd_pr__pfet_01v8_J8PPQP  XM9
timestamp 1755446217
transform 1 0 3927 0 1 -8107
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_X8MKUN  XM10
timestamp 1755446217
transform 1 0 2457 0 1 -8165
box -263 -269 263 269
use sky130_fd_pr__nfet_01v8_TGNW9T  XM11
timestamp 1755446217
transform 1 0 4615 0 1 -8762
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_J8PPQP  XM12
timestamp 1755446217
transform 1 0 4929 0 1 -8105
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_TGNW9T  XM13
timestamp 1755446217
transform 1 0 4931 0 1 -8762
box -211 -310 211 310
<< labels >>
flabel metal1 5154 -7852 5354 -7652 0 FreeSans 256 0 0 0 OUT
port 2 nsew
rlabel metal1 5212 -9170 5412 -8970 1 VSS
port 4 n
rlabel metal1 3118 -7836 3318 -7636 1 VDD
port 3 n
flabel metal1 2312 -9176 2512 -8976 0 FreeSans 256 0 0 0 IN1
port 0 nsew
flabel metal1 2730 -9176 2930 -8976 0 FreeSans 256 0 0 0 IN2
port 1 nsew
<< end >>
