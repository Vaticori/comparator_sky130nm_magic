magic
tech sky130A
timestamp 1753299038
<< error_p >>
rect -2 4 4 29
rect -27 -2 -2 4
rect 4 -2 29 4
rect -2 -27 4 -2
<< varactor >>
rect -2 -2 4 4
<< end >>
