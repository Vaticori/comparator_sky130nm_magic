magic
tech sky130A
magscale 1 2
timestamp 1754957036
<< error_s >>
rect 3848 -7830 4006 -7824
rect 3848 -7850 3854 -7830
rect 4000 -7850 4006 -7830
rect 3848 -7856 4006 -7850
<< pwell >>
rect 1940 -8608 2006 -8556
rect 2256 -8608 2322 -8556
rect 2572 -8610 2638 -8560
rect 2888 -8608 2954 -8556
rect 3470 -8620 3536 -8562
rect 3312 -8660 3376 -8644
rect 3624 -8650 3706 -8634
rect 2668 -8800 2864 -8678
rect 3312 -8838 3476 -8660
rect 3624 -8662 3796 -8650
rect 3312 -8866 3376 -8838
rect 3530 -8842 3796 -8662
rect 3624 -8844 3796 -8842
rect 3624 -8860 3706 -8844
rect 3920 -8846 3934 -8606
rect 3952 -8662 4006 -8646
rect 3952 -8844 4108 -8662
rect 3952 -8856 4008 -8844
rect 2698 -8922 2828 -8906
rect 3470 -8940 3538 -8880
rect 3786 -8938 3854 -8878
rect 4100 -8938 4168 -8878
rect 2698 -9088 2828 -9066
rect 3404 -9082 3596 -8968
rect 4696 -9038 4706 -8994
rect 4846 -9038 4872 -8986
rect 4220 -9108 5046 -9038
<< locali >>
rect 4436 -8072 4472 -7918
rect 3328 -8838 3362 -8660
rect 4442 -8672 4474 -8584
rect 4442 -8940 4474 -8858
<< viali >>
rect 3848 -7856 4006 -7824
rect 4534 -7856 5008 -7820
rect 3752 -8196 3786 -8018
rect 4436 -8290 4472 -8072
rect 2114 -8794 2148 -8700
rect 2746 -8790 2780 -8692
rect 3642 -8842 3680 -8648
rect 3960 -8838 3994 -8662
rect 4442 -8858 4476 -8672
rect 3422 -9024 3582 -8990
rect 3740 -9024 3900 -8990
rect 4054 -9026 4214 -8992
rect 4536 -9036 4696 -9002
rect 4852 -9036 5010 -9002
<< metal1 >>
rect 4518 -7722 5018 -7720
rect 2392 -7780 5018 -7722
rect 3770 -7788 5018 -7780
rect 4518 -7820 5018 -7788
rect 4518 -7856 4534 -7820
rect 5008 -7856 5018 -7820
rect 4518 -7872 5018 -7856
rect 1934 -7912 2652 -7908
rect 1934 -7962 2970 -7912
rect 3578 -7976 3644 -7910
rect 3894 -7976 3960 -7910
rect 4352 -7974 4646 -7908
rect 4686 -7974 4960 -7908
rect 3732 -8018 3902 -8008
rect 3732 -8196 3752 -8018
rect 3786 -8196 3902 -8018
rect 4352 -8020 4392 -7974
rect 4426 -7976 4488 -7974
rect 4686 -7978 4788 -7974
rect 4686 -8002 4724 -7978
rect 3952 -8072 4392 -8020
rect 4426 -8070 4492 -8060
rect 4534 -8070 4592 -8006
rect 4426 -8072 4592 -8070
rect 3732 -8210 3902 -8196
rect 1932 -8288 2968 -8238
rect 3578 -8304 3644 -8238
rect 3894 -8304 3960 -8238
rect 4164 -8432 4236 -8072
rect 4426 -8290 4436 -8072
rect 4472 -8208 4592 -8072
rect 4640 -8206 4724 -8002
rect 4472 -8290 4484 -8208
rect 4894 -8240 4962 -8236
rect 4426 -8306 4484 -8290
rect 3892 -8470 4238 -8432
rect 1940 -8608 2006 -8556
rect 2256 -8608 2322 -8556
rect 2572 -8610 2638 -8554
rect 2888 -8608 2954 -8556
rect 3470 -8620 3536 -8562
rect 3786 -8620 3852 -8562
rect 3892 -8606 3934 -8470
rect 1998 -8690 2046 -8640
rect 2216 -8690 2262 -8640
rect 3624 -8648 3706 -8634
rect 1998 -8700 2262 -8690
rect 1998 -8794 2114 -8700
rect 2148 -8794 2262 -8700
rect 1998 -8800 2262 -8794
rect 2668 -8692 2864 -8678
rect 2668 -8790 2746 -8692
rect 2780 -8790 2864 -8692
rect 2668 -8800 2864 -8790
rect 1998 -8840 2046 -8800
rect 2216 -8840 2262 -8800
rect 3430 -8838 3476 -8660
rect 3624 -8662 3642 -8648
rect 3530 -8842 3642 -8662
rect 3680 -8650 3706 -8648
rect 3892 -8650 3920 -8606
rect 4102 -8620 4168 -8562
rect 4582 -8576 4646 -8246
rect 4894 -8306 4964 -8240
rect 4896 -8574 4964 -8306
rect 5842 -8546 6042 -8346
rect 4582 -8632 4650 -8576
rect 4686 -8632 4964 -8574
rect 4686 -8634 4924 -8632
rect 3680 -8842 3796 -8650
rect 3874 -8652 3920 -8650
rect 3624 -8844 3796 -8842
rect 3624 -8860 3706 -8844
rect 3844 -8846 3920 -8652
rect 3952 -8662 4006 -8646
rect 4686 -8656 4722 -8634
rect 3952 -8838 3960 -8662
rect 3994 -8838 4108 -8662
rect 3952 -8844 4108 -8838
rect 4432 -8672 4488 -8656
rect 3952 -8856 4006 -8844
rect 4432 -8858 4442 -8672
rect 4476 -8674 4488 -8672
rect 4676 -8674 4722 -8656
rect 4476 -8856 4590 -8674
rect 4642 -8850 4722 -8674
rect 4476 -8858 4488 -8856
rect 1918 -8920 2954 -8870
rect 2082 -9066 2174 -8920
rect 2698 -8922 2828 -8920
rect 2710 -9066 2820 -8922
rect 3470 -8940 3538 -8880
rect 3786 -8938 3854 -8878
rect 4100 -8938 4168 -8878
rect 4432 -8882 4488 -8858
rect 4582 -8946 4650 -8890
rect 4896 -8948 4964 -8892
rect 3404 -8990 3596 -8968
rect 3404 -9024 3422 -8990
rect 3582 -9024 3596 -8990
rect 3404 -9040 3596 -9024
rect 3722 -8990 3914 -8970
rect 3722 -9024 3740 -8990
rect 3900 -9024 3914 -8990
rect 3722 -9040 3914 -9024
rect 4036 -8992 4228 -8970
rect 4036 -9026 4054 -8992
rect 4214 -9026 4228 -8992
rect 4036 -9038 4228 -9026
rect 4526 -9002 4706 -8986
rect 4526 -9036 4536 -9002
rect 4696 -9036 4706 -9002
rect 4846 -9002 5022 -8986
rect 4846 -9036 4852 -9002
rect 5010 -9036 5022 -9002
rect 4526 -9038 5022 -9036
rect 4036 -9040 5046 -9038
rect 2032 -9266 2232 -9066
rect 2662 -9266 2862 -9066
rect 3402 -9108 5046 -9040
rect 3402 -9110 4228 -9108
<< metal2 >>
rect 3452 -8620 4184 -8570
use 1meg  R2
timestamp 0
transform 1 0 4744 0 1 -8517
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_V8CAV6  sky130_fd_pr__nfet_01v8_V8CAV6_0
timestamp 1754957036
transform 1 0 2605 0 1 -8740
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  sky130_fd_pr__nfet_01v8_V8CAV6_1
timestamp 1754957036
transform 1 0 1973 0 1 -8740
box -211 -310 211 310
use sky130_fd_pr__cap_mim_m3_1_3E28FE  XC8
timestamp 1754957036
transform 0 -1 5494 1 0 -8436
box -686 -240 686 240
use sky130_fd_pr__nfet_01v8_V8CAV6  XM1
timestamp 1754957036
transform 1 0 3503 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XM2
timestamp 1754957036
transform 1 0 2921 0 1 -8740
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM3
timestamp 1754957036
transform 1 0 3611 0 1 -8107
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM4
timestamp 1754957036
transform 1 0 4613 0 1 -8105
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_V8CAV6  XM5
timestamp 1754957036
transform 1 0 4135 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM6
timestamp 1754957036
transform 1 0 2605 0 1 -8101
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_V8CAV6  XM7
timestamp 1754957036
transform 1 0 3819 0 1 -8750
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XM8
timestamp 1754957036
transform 1 0 2289 0 1 -8740
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM9
timestamp 1754957036
transform 1 0 3927 0 1 -8107
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM10
timestamp 1754957036
transform 1 0 2921 0 1 -8101
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_V8CAV6  XM11
timestamp 1754957036
transform 1 0 4615 0 1 -8762
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XUW9MZ  XM12
timestamp 1754957036
transform 1 0 4929 0 1 -8105
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_V8CAV6  XM13
timestamp 1754957036
transform 1 0 4931 0 1 -8762
box -211 -310 211 310
<< labels >>
flabel metal1 2032 -9266 2232 -9066 0 FreeSans 256 0 0 0 IN1
port 0 nsew
flabel metal1 5842 -8546 6042 -8346 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 2662 -9266 2862 -9066 0 FreeSans 256 0 0 0 IN2
port 1 nsew
<< end >>
